module RISCV_tb();
reg clk;
reg rst;

parameter CLK_PERIOD=20;
riscv DUT(
.clk(clk),
.rst(rst)
);

initial
begin
forever
#(CLK_PERIOD/2) clk=~clk;
end
initial 
begin
clk=1'b0;
rst=1'b0;
#(CLK_PERIOD);
rst=1'b1;
#(CLK_PERIOD);
#1000;
$finish;
end
endmodule
