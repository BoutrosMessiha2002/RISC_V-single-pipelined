module ALU #( parameter DATA=32, parameter CONTROL=3)(
input [DATA-1:0] SrcA,
input [DATA-1:0] SrcB,
input [CONTROL-1:0] ALUControl,
output reg [DATA-1:0] ALUResult,
output zero
);

always @(*)
begin
case (ALUControl)
3'b000: ALUResult=SrcA+SrcB;
3'b001: ALUResult=SrcA-SrcB;
3'b010: ALUResult=SrcA&SrcB;
3'b011: ALUResult=SrcA|SrcB;
3'b101: ALUResult=SrcA<SrcB;
default: ALUResult='b0;
endcase
end
assign zero=((SrcA-SrcB)=='b0);
endmodule
