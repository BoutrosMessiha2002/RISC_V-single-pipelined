module riscv(
input clk,
input rst
);
wire [31:0] PCNext;
wire [31:0] PC;
wire [31:0] Instr;
wire [31:0] PCPlus4;
wire [31:0] SrcA;
wire [31:0] SrcB;
wire [31:0] ALUResult;
wire [31:0] ReadData;
wire [31:0] Result;
wire [31:0] ImmExt;
wire [31:0] PCTarget;
wire [31:0] WriteData;
wire PCSrc;
wire [1:0] ResultSrc;
wire MemWrite;
wire [2:0] ALUControl;
wire ALUSrc;
wire [1:0] ImmSrc;
wire RegWrite;
wire zero;
mux2to1 #(.DATA(32))PCmux(
.A(PCPlus4),
.B(PCTarget),
.sel(PCSrc),
.out(PCNext)
);

PC PC_dut(
.clk(clk),
.rst(rst),
.PC(PC),
.PCNext(PCNext)
);

adder adder_4(
.A(PC),
.B(32'd4),
.out(PCPlus4)
);

instr_mem #(.ADDRESS(32), .INSTR(32))instr_m(
.A(PC),
.RD(Instr)
);

reg_file#(.ADDRESS(5), .DATA(32)) reg_f(
.clk(clk),
.A1(Instr[19:15]),
.A2(Instr[24:20]),
.A3(Instr[11:7]),
.WD3(Result),
.WE3(RegWrite),
.RD1(SrcA),
.RD2(WriteData)
);

mux2to1 #(.DATA(32))SrcB_mux(
.A(WriteData),
.B(ImmExt),
.sel(ALUSrc),
.out(SrcB)
);

sign_extend ext(
.in_val(Instr[31:7]),
.ImmExt(ImmExt),
.ImmSrc(ImmSrc)
);

adder adder_ext(
.A(PC),
.B(ImmExt),
.out(PCTarget)
);

ALU #(.DATA(32), .CONTROL(3))ALU_dut(
.SrcA(SrcA),
.SrcB(SrcB),
.zero(zero),
.ALUResult(ALUResult),
.ALUControl(ALUControl)
);

data_mem #(.ADDRESS(128),.DATA(32), .N(128))data(
.A(ALUResult),
.WD(WriteData),
.clk(clk),
.WE(MemWrite),
.RD(ReadData)
);

 mux4to1 #(.DATA(32)) read_mux(
.A(ALUResult),
.B(ReadData),
.C(PCPlus4),
.sel(ResultSrc),
.out(Result)
);

control_unit control(
.op(Instr[6:0]),
.funct3(Instr[14:12]),
.funct7_5(Instr[30]),
.zero(zero),
.PCSrc(PCSrc),
.ResultSrc(ResultSrc),
.MemWrite(MemWrite),
.ALUControl(ALUControl),
.ALUSrc(ALUSrc),
.ImmSrc(ImmSrc),
.RegWrite(RegWrite)
);
endmodule


